li x10 10
li x11 10
nop
nop
nop
nop
nop
beq x10 x11 label
li x12 33
li x13 33
label:
li x14 33
li x15 33