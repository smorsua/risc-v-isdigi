`ifndef OPERATION_TYPE_HEADER
`define OPERATION_TYPE_HEADER
enum bit [3:0] { ADD, SLT, SLTU, AND, OR, XOR, LUI, AUIPC, SUB, BEQ, BNE,
LW, SW } e_operations;
`endif OPERATION_TYPE_HEADER