`ifndef OPERATION_TYPE_HEADER
`define OPERATION_TYPE_HEADER
typedef enum { 
	ADD, 
	SUB, 
	LESS_THAN, 
	GREATER_OR_EQUAL_THAN, 
	AND,
	OR, 
	XOR, 
	LEFT_SHIFT, 
	SIGNED_LEFT_SHIFT, 
	RIGHT_SHIFT, 
	SIGNED_RIGHT_SHIFT } e_operations;
`endif OPERATION_TYPE_HEADER