module CONTROL(
    input [6:0] INSTRUCTION_FORMAT,
    output BRANCH,
    output MEM_READ,
    output MEM_TO_REG,
    output ALU_OP,
    output MEM_WRITE,
    output ALU_SRC,
    output REG_WRITE
);
endmodule