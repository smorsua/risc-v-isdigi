module ALU_CONTROL(
    input [3:0] funct3And30
    input ALUOp,
    output [3.0] ALUSelection
);


    

endmodule 