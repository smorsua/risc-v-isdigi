`ifndef OPERATION_TYPE_HEADER
`define OPERATION_TYPE_HEADER
enum bit [3:0] { ADD, SUB, LESS_THAN, GREATER_OR_EQUAL_THAN, AND, OR, XOR, LEFT_SHIFT, RIGHT_SHIFT } e_operations;
`endif OPERATION_TYPE_HEADER